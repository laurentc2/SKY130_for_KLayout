* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.SUBCKT sky130_fd_sc_hs__and2_1 A B VGND VNB VPWR VPB X
*.PININFO A:I B:I VGND:I VNB:I VPB:I VPWR:I X:O
MMP0 y A VPWR VPB pfet_01v8 w=0.84 l=0.15
MMP1 y B VPWR VPB pfet_01v8 w=0.84 l=0.15
MMIP0 X y VPWR VPB pfet_01v8 w=1.12 l=0.15
MMN0 y A sndA VNB nfet_01v8_lvt w=0.64 l=0.15
MMN1 sndA B VGND VNB nfet_01v8_lvt w=0.64 l=0.15
MMIN0 X y VGND VNB nfet_01v8_lvt w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__and2_1


.SUBCKT sky130_fd_sc_hs__and2_2 A B VGND VNB VPWR VPB X
*.PININFO A:I B:I VGND:I VNB:I VPB:I VPWR:I X:O
MMP0 y A VPWR VPB pfet_01v8 w=1.0 l=0.15
MMP1 y B VPWR VPB pfet_01v8 w=1.0 l=0.15
MMIP0 X y VPWR VPB pfet_01v8 m=2 w=1.12 l=0.15
MMN0 y A sndA VNB nfet_01v8_lvt w=0.74 l=0.15
MMN1 sndA B VGND VNB nfet_01v8_lvt w=0.74 l=0.15
MMIN0 X y VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__and2_2


.SUBCKT sky130_fd_sc_hs__and2_4 A B VGND VNB VPWR VPB X
*.PININFO A:I B:I VGND:I VNB:I VPB:I VPWR:I X:O
MMP0 y A VPWR VPB pfet_01v8 m=2 w=0.84 l=0.15
MMP1 y B VPWR VPB pfet_01v8 m=2 w=0.84 l=0.15
MMIP0 X y VPWR VPB pfet_01v8 m=4 w=1.12 l=0.15
MMN0 y A sndA VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMN1 sndA B VGND VNB nfet_01v8_lvt m=2 w=0.64 l=0.15
MMIN0 X y VGND VNB nfet_01v8_lvt m=4 w=0.74 l=0.15
.ENDS sky130_fd_sc_hs__and2_4
